------------------------------------------------------------------------------------
---- Company: nope
---- Engineer: me
---- 
---- Create Date:    13:48:22 10/06/2016 
---- Design Name: 
---- Module Name:    cleaner - Behavioral 
---- Project Name: 
---- Target Devices: 
---- Tool versions: 
---- Description: 
----
---- Dependencies: 
----
---- Revision: 
---- Revision 0.01 - File Created
---- Additional Comments: 
----
------------------------------------------------------------------------------------
--
----type servo_in_type is record
----    pos_i : std_logic_vector(10 downto 0);
----end record;
----
----type servo_out_type is record
----    servo_o : std_logic;
----end record;
--library IEEE;
--use IEEE.STD_LOGIC_1164.all;
--
--
--package servo_comp is
--
--component servo is
--  Port ( clk_i : in  STD_LOGIC;
--         reset_i : in STD_LOGIC;
--         pos_i : in std_logic_vector(10 downto 0);
--         servo_o : out std_logic
--         );
--end component;
--
--end package;
--
--
--library IEEE;
--use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.STD_LOGIC_UNSIGNED.ALL;
--use IEEE.NUMERIC_STD.ALL;
--
--library UNISIM;
--use UNISIM.VComponents.all;
--
--entity servo is
--  Port ( clk_i : in  STD_LOGIC;
--         reset_i : in STD_LOGIC;
--         pos_i : in std_logic_vector(10 downto 0);
--         servo_o : out std_logic);
--end servo;
--
----------------------------------------------------------------------------------
----------------------------------------------------------------------------------
--architecture twoproc of servo is
--
--  signal clk_1MHz : std_logic;
--  constant REPETITIONS: integer := 30000;
--  constant T20MS: integer := 20_000;
--  --signal pos_i : std_logic_vector(10 downto 0) := std_logic_vector(to_unsigned(1000,11));
--  signal cnt : std_logic_vector(10 downto 0) := "00000000000";
--  signal counting : std_logic;
--  signal h : std_logic;
--  signal d2 : std_logic;
--  signal d3 : std_logic;
--  signal reported : std_logic_vector(10 downto 0);
--
--begin
--
------------------------------------------------------------------------------------
---- Digital Clock Manager
----
---- sensitivity : clk_i
---- extra inputs:
---- outputs     : clk_1MHz
------------------------------------------------------------------------------------
--  DCM_SP_1MHz : DCM_SP
--    generic map (
--      CLKFX_DIVIDE   => 24, 
--      CLKFX_MULTIPLY => 2
--      )
--    port map (
--      CLKFX => clk_1MHz,  --  1MHz out
--      CLKIN => clk_i,     -- 12MHz in
--      RST   => reset_i
--      );
--
--
--
--  comb : process(reset_i, pos_i, clk_1MHz) is
--    variable counter : integer := 0;
--    variable rep : integer := REPETITIONS;
--  begin
--    if reset_i = '1' then
--      rep := REPETITIONS;
--      counter := 0;
--      servo_o <= '0';
--      h <= '0';
--    else
--      if rising_edge(clk_1MHz) then
--        if counter = T20MS then -- 50Hz trigger
--          if rep > 0 then
--            rep := rep - 1;
--            servo_o <= '1';
--            h <= '1';
--          end if;
--          counter := 0;
--        end if;
--        if counter = pos_i then
--          servo_o <= '0';
--          h <= '0';
--        end if;
--        counter := counter + 1;
--      elsif falling_edge(clk_1MHz) then
--        -- do nothing;
--      else --pos_i changed
--        rep := REPETITIONS;
--      end if;
--    end if;
--  end process;
--
--
--------------------------------------------------------------------------------------
------ DIJON pulse measurement
------
------ sensitivity : servo_helper, clk_1MHz, reset_i
------ extra inputs: 
------ outputs     : p1, p2
--------------------------------------------------------------------------------------  
--
--test_counter_a_pw: process(clk_1Mhz) -- Synchronous process depends ONLY on clock edge
--begin
--  if clk_1MHz'event and clk_1MHz='1' then -- Synchronous process, clock edge is outer "if"
--      d2 <= h;  -- First D FF stage (common synchronization point)
--      d3 <= d2; -- Second D FF stage for edge detect
--      if  d3 = '0' and d2 = '1' then -- Detect rising edge
--        cnt <= "00000000000";
--      elsif d3 = '1' and d2 = '0' then -- Detect falling edge
--        reported <= cnt + 1;  -- Capture count
--      else
--        cnt <= cnt + 1;
--      end if;
--    end if;
--end process test_counter_a_pw;
--
--
--end twoproc;
